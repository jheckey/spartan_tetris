
module scanline_fifo (
    input   wire        clk,
    input   wire        rst,
    input   wire        din,
    input   reg  [23:0] pixin,
    output  reg  [2:0]  pixout
);

reg     [23:0]  buffer;


endmodule

