
module siggen (
    input   wire        clk,        // 50MHz
    input   wire        rst,
    input   wire [10:0] cnt_X,
    input   wire [9:0]  cnt_Y,
    output  reg  [47:0] pixels
);

localparam XOFFSET = 8;		// 224 clks before visible pixels; 224/(16 pix/tile * 2 clks/pix) = 7; +1 to start before the tile needed
localparam YOFFSET = 12;	// 12 lines scanned above display area

// 640 / 16 = 40
// 480 / 16 = 30
wire	  [9:0]   offset_y = cnt_Y - YOFFSET;		// Reset to start of display area
wire    [5:0]   tile_x 	 = cnt_X[10:5] - XOFFSET;
wire    [5:0]   tile_y 	 = offset_y[9:4];
reg     [47:0]  pixels_n;

always @(posedge clk or posedge rst) begin
    if (rst) begin
        pixels  <= 48'd0;
    end
    else begin
        pixels  <= pixels_n;
    end
end

always @* begin
	pixels_n = {8{{tile_y[2:0],tile_x[2:0]}}};
	/*
	case (tile_y)
		0:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		1:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		2:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		3:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		4:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		5:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		6:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		7:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		8:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		9:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		10:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		11:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		12:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		13:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		14:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		15:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		16:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		17:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		18:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		19:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		20:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		21:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		22:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		23:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		24:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		25:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		26:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		27:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		28:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		29:
			case (tile_x)
				0:  pixels_n = {16{3'b001}};
				1:  pixels_n = {16{3'b010}};
				2:  pixels_n = {16{3'b100}};
				3:  pixels_n = {16{3'b001}};
				4:  pixels_n = {16{3'b010}};
				5:  pixels_n = {16{3'b100}};
				6:  pixels_n = {16{3'b001}};
				7:  pixels_n = {16{3'b010}};
				8:  pixels_n = {16{3'b100}};
				9:  pixels_n = {16{3'b001}};
				10:  pixels_n = {16{3'b010}};
				11:  pixels_n = {16{3'b100}};
				12:  pixels_n = {16{3'b001}};
				13:  pixels_n = {16{3'b010}};
				14:  pixels_n = {16{3'b100}};
				15:  pixels_n = {16{3'b001}};
				16:  pixels_n = {16{3'b010}};
				17:  pixels_n = {16{3'b100}};
				18:  pixels_n = {16{3'b001}};
				19:  pixels_n = {16{3'b010}};
				20:  pixels_n = {16{3'b100}};
				21:  pixels_n = {16{3'b001}};
				22:  pixels_n = {16{3'b010}};
				23:  pixels_n = {16{3'b100}};
				24:  pixels_n = {16{3'b001}};
				25:  pixels_n = {16{3'b010}};
				26:  pixels_n = {16{3'b100}};
				27:  pixels_n = {16{3'b001}};
				28:  pixels_n = {16{3'b010}};
				29:  pixels_n = {16{3'b100}};
				30:  pixels_n = {16{3'b001}};
				31:  pixels_n = {16{3'b010}};
				32:  pixels_n = {16{3'b100}};
				33:  pixels_n = {16{3'b001}};
				34:  pixels_n = {16{3'b010}};
				35:  pixels_n = {16{3'b100}};
				36:  pixels_n = {16{3'b001}};
				37:  pixels_n = {16{3'b010}};
				38:  pixels_n = {16{3'b100}};
				39:  pixels_n = {16{3'b001}};
			endcase
		default: pixels_n = {16{3'b101}};
	endcase
	*/
end

endmodule

